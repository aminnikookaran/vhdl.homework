module Simple_Dual_Port_Ram_1024x8bit_Ent (iwA,iadrA,iclkA,idataA,irB,iadrB,iclkB,odataB);
input iwA;
input [9:0]iadrA;
input iclkA;
input [7:0]idataA;
input irB;
input [9:0]iadrB;
input iclkB;
output [7:0]odataB;
endmodule

